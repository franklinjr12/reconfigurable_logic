library verilog;
use verilog.vl_types.all;
entity vhdl_test_vlg_check_tst is
    port(
        C               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end vhdl_test_vlg_check_tst;
