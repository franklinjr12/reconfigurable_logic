library verilog;
use verilog.vl_types.all;
entity calcula_seno_vlg_vec_tst is
end calcula_seno_vlg_vec_tst;
