library verilog;
use verilog.vl_types.all;
entity vhdl_test is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : out    vl_logic
    );
end vhdl_test;
