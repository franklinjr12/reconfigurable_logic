library verilog;
use verilog.vl_types.all;
entity vhdl_test_vlg_vec_tst is
end vhdl_test_vlg_vec_tst;
