library verilog;
use verilog.vl_types.all;
entity my_jk_vlg_vec_tst is
end my_jk_vlg_vec_tst;
